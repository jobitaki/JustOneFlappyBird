`default_nettype none

module uniprocessor();

endmodule: uniprocessor